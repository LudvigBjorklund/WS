library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.num_of_bits.all;


package DT_IDs is


end package DT_IDs;



