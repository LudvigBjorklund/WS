
-- -- Import necessary libraries
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Include the Altera megafunction components library
-- For Synthesis, ensure the Altera libraries are available in your project settings
-- library altera_mf;
-- use altera_mf.altera_mf_components.all;

entity tbl_read_ow_sim is 
    generic(
        table_name : string := "R0";
        hex_init : string := "LUT_2D.hex"  -- Name of the HEX (or MIF) file for initialization
    );
    port(
        i_clk   : in  std_logic;                     -- Clock signal
        i_raddr : in  unsigned(7 downto 0);            -- Read address (8-bit)
        i_waddr : in  unsigned(7 downto 0);            -- Write address (8-bit)
        i_wr_en : in  std_logic;                        -- Write enable signal
        i_data  : in  unsigned(15 downto 0);           -- 16-bit data input for writez
        o_data  : out unsigned(15 downto 0)            -- 16-bit data output for read
    );
end entity tbl_read_ow_sim;

architecture rtl of tbl_read_ow_sim is
    -- Internal signal to connect the megafunction's output
    signal mem_out : std_logic_vector(15 downto 0);



type flat_lut is array (0 to 175) of unsigned(15 downto 0);

signal r_R0tbl : flat_lut := (
  -- Row 0 (Address 0 to 10)
  "0111111100000000", "0011001000000000", "0010001100000000", "0001100100000000", "0001000100000000", "0000111100000000", "0000111000000000", "0000110100000000", "0000110010000000", "0000101100000000", "0000100100000000",
  -- Row 1 (Address 11 to 21)
  "0111110100000000", "0010100000000000", "0001101100000000", "0001010000000000", "0001000000000000", "0000111000000000", "0000110000000000", "0000101100000000", "0000101000000000", "0000100100000000", "0000100000000000",
  -- Row 2 (Address 22 to 32)
  "0111101100000000", "0010000000000000", "0001100000000000", "0001001100000000", "0000111100000000", "0000110100000000", "0000101100000000", "0000101000000000", "0000100110000000", "0000100010000000", "0000011110000000",
  -- Row 3
  "0111100000000000", "0001100100000000", "0001011000000000", "0001001000000000", "0000111000000000", "0000110000000000", "0000101010000000", "0000100110000000", "0000100010000000", "0000011100000000", "0000011000000000",
  -- Row 4
  "0110111000000000", "0001010000000000", "0001001000000000", "0001000100000000", "0000110100000000", "0000101100000000", "0000101000000000", "0000100100000000", "0000011111000000", "0000011011000000", "0000010110000000",
  -- Row 5
  "0101111100000000", "0001000100000000", "0000111100000000", "0000111000000000", "0000110000000000", "0000101000000000", "0000100100000000", "0000100000000000", "0000011101000000", "0000011010000000", "0000010101000000",
  -- Row 6
  "0101000000000000", "0001000000000000", "0000111000000000", "0000110100000000", "0000101100000000", "0000100100000000", "0000100000000000", "0000011110000000", "0000011100000000", "0000011001000000", "0000010100100000",
  -- Row 7
  "0100011100000000", "0000111100000000", "0000110100000000", "0000110000000000", "0000101000000000", "0000011110000000", "0000011011000000", "0000011010000000", "0000011001000000", "0000011000000000", "0000010100000000",
  -- Row 8
  "0011111100000000", "0000111000000000", "0000110000000000", "0000101000000000", "0000100101000000", "0000011000000000", "0000010111000000", "0000010110000000", "0000010101100000", "0000010100100000", "0000010011100110",
  -- Row 9
  "0011011000000000", "0000110100000000", "0000101100000000", "0000100110000000", "0000100100000000", "0000010100000000", "0000010011000000", "0000010010000000", "0000010001000000", "0000010000100000", "0000010000000000",
  -- Row 10
  "0010111100000000", "0000110010000000", "0000101010000000", "0000100100000000", "0000100000000000", "0000010010000000", "0000010001100000", "0000010001000000", "0000010000100110", "0000010000000000", "0000001111100000",
  -- Row 11
  "0010100100000000", "0000110000000000", "0000101000000000", "0000100000000000", "0000011100000000", "0000010000000000", "0000001111100000", "0000001111000000", "0000001110100000", "0000001110000000", "0000001101100110",
  -- Row 12
  "0010010000000000", "0000101100000000", "0000100110000000", "0000011110000000", "0000011000000000", "0000001111000000", "0000001110000000", "0000001101100000", "0000001100100000", "0000001100000000", "0000001011100110",
  -- Row 13
  "0010000100000000", "0000101000000000", "0000100100000000", "0000011100000000", "0000010110000000", "0000001101000000", "0000001100100000", "0000001100000000", "0000001011100110", "0000001011100001", "0000001011001100",
  -- Row 14
  "0001111000000000", "0000100100000000", "0000100010000000", "0000011010000000", "0000010100000000", "0000001100000000", "0000001011001100", "0000001011000000", "0000001010110011", "0000001010101011", "0000001010011001",
  -- Row 15
  "0001110000000000", "0000011100000000", "0000011011001100", "0000011001001100", "0000010011100110", "0000001011000000", "0000001010011001", "0000001010001100", "0000001010000000", "0000001001110011", "0000001001100110"
);


signal r_a1 :flat_lut := (
  -- Row 0
  "0001100111011010", "0010100011110101", "0101000111101011", "0101000011101000", "0110001110101000", "0110100110110100", "0111000111000111", "0110101100010101", "0110001101001100", "0101110100010111", "0100101001001101",
  -- Row 1
  "0001110101110110", "0010011001111110", "0100110011111100", "0100110111000011", "0011111000101010", "0011110001110010", "0100100001011110", "0101001001011111", "0100110011011100", "0011100110001100", "0011100011100111",
  -- Row 2
  "0001111011001100", "0010001100001000", "0101000011010111", "0101011110010100", "0010010001011010", "0011100101111100", "0100001100000000", "0101001001111010", "0100110000000100", "0011101001000011", "0011100000100111",
  -- Row 3
  "0001011110111110", "0010101000010111", "0110000001110110", "0100100101111111", "0010010101111000", "0011100000111001", "0011111011100000", "0101001000000101", "0100101101110100", "0011101000011001", "0011011111100100",
  -- Row 4
  "0001010110101100", "0011001010110110", "0111100010111110", "0100011001101111", "0010011001110100", "0011011101011001", "0011111001111010", "0101000101100110", "0100101101010100", "0011101001000011", "0011100000111010",
  -- Row 5
  "0001110000111111", "0100010011011010", "0111001011000010", "0100100000000001", "0010011100111001", "0011011100111111", "0011111001011000", "0101000100111110", "0100101000000110", "0011101000100101", "0011011111100001",
  -- Row 6
  "0010001001011001", "0100010101001001", "0110101110100100", "0100101111010011", "0010100000101101", "0011011110000000", "0011110111011011", "0101000011010001", "0100100110001101", "0011101000001100", "0011011101001101",
  -- Row 7
  "0010100000101000", "0100100111110100", "0110100000000000", "0101000010101101", "0010100110011010", "0011011011110110", "0011110111001111", "0100111111111101", "0100100000111110", "0011100101011101", "0011011010111000",
  -- Row 8
  "0010111010001011", "0100100010011100", "0110101011000111", "0101010011101100", "0010101000101111", "0011010110101010", "0011110001010100", "0100110110010001", "0100011110111000", "0011101010010001", "0011011111010000",
  -- Row 9
  "0011011010011101", "0100001010001111", "0110010100110110", "0100110000010110", "0010011110010001", "0011011100010010", "0011111000010100", "0101001001110110", "0100100111101111", "0011110101110110", "0011110100110001",
  -- Row 10
  "0011100011100011", "0011111101100011", "0101110101011011", "0100101100111010", "0010011110000011", "0011100101100101", "0100000101001000", "0101001101110001", "0100101100111001", "0100010011110100", "0100000010101001",
  -- Row 11
  "0100000001111010", "0101011001110001", "0101101111001001", "0100110010010010", "0010011110110001", "0100000000000000", "0100100101100111", "0101100100111100", "0100111100001110", "0101000000000000", "0100110001111101",
  -- Row 12
  "0100101111011010", "0110101001111110", "0101111011111010", "0100110101011001", "0010100001010000", "0100111000000100", "0101011011111010", "0110100111101000", "0101111010010001", "0110000110000110", "0101111111100000",
  -- Row 13
  "0101000000101000", "0111001101000001", "0110001011011001", "0100111111111001", "0010100100111100", "0110000110000110", "0110101110010111", "0111111101111011", "0111011000110101", "0111100111100111", "0111010111110001",
  -- Row 14
  "0101000011101000", "0111110010001110", "0110000010010110", "0011111100110010", "0010111111000100", "0011010101010101", "0100010011110100", "0100000011000100", "0011111110100110", "0011111100110101", "0011110111101011",
  -- Row 15
  "0100110100011001", "1000110111111110", "0110110100111010", "0011100011100011", "0011010000000011", "0100011100111100", "0101001010111111", "0101000001010000", "0101000000010100", "0101110100010100", "0101110001110111"
);
signal r_c1 : flat_lut := (
 -- Row 0 
 "0100111011000100", "0100000000000000", "0011001100110011", "0010010111101101", "0010010101011111", "0010000100001000", "0010000000000000", "0001110001110001", "0001100110011001", "0001011101000101", "0001001001001001",
 -- Row 1 
 "0100110001101010", "0011001100110011", "0010100011110101", "0001111100000111", "0001001111011000", "0001001001101010", "0001001111011000", "0001010101010101", "0001001101010010", "0000111000000111", "0000110110100111",
 -- Row 2 
 "0100100100100100", "0010101010101010", "0010011101100010", "0010000000000000", "0001001011110110", "0001000100010001", "0001000111100110", "0001010011010000", "0001001010011110", "0000110111010110", "0000110100100000",
 -- Row 3 
 "0011001100110011", "0010111010001011", "0010101010101010", "0001100001100001", "0001001001001001", "0001000010000100", "0001000010011111", "0001010001111010", "0001001001001001", "0000110110100111", "0000110011101101",
 -- Row 4 
 "0010101010101010", "0011001100110011", "0011000011000011", "0001010101010101", "0001000110100111", "0001000000000000", "0001000001000001", "0001010000000000", "0001000111110111", "0000110101111001", "0000110011001100",
 -- Row 5 
 "0011001100110011", "0100000000000000", "0010101010101010", "0001010000010100", "0001000100010001", "0000111111000000", "0001000000000000", "0001001110110001", "0001000101101010", "0000110101000011", "0000110010001100",
 -- Row 6 
 "0011100011100011", "0011101011011001", "0010010010010010", "0001001101010010", "0001000010000100", "0000111110011100", "0000111110101000", "0001001101010010", "0001000100010001", "0000110100001111", "0000110000111111",
 -- Row 7 
 "0011110000111100", "0011100011100011", "0010000000000000", "0001001010011110", "0001000000011001", "0000111101010100", "0000111110000011", "0001001011110110", "0001000010011111", "0000110011001100", "0000110000000100",
 -- Row 8 
 "0100000000000000", "0011001100110011", "0001111000011110", "0001000111110111", "0000111110000011", "0000111011100010", "0000111100001111", "0001001001001001", "0001000001101001", "0000110011111110", "0000110000110000",
 -- Row 9 
 "0100010001000100", "0010101010101010", "0001110101000001", "0001000100111101", "0000111100100101", "0000111010100000", "0000111011010111", "0001001010011110", "0001000000110011", "0000110100001111", "0000110011001100",
 -- Row 10 
 "0100000000000000", "0010010010010010", "0001110001110001", "0001000111110111", "0000111110011100", "0000111011001100", "0000111100100101", "0001001001001001", "0001000000000000", "0000111000111000", "0000110100100000",
 -- Row 11 
 "0100001001111110", "0010110110110110", "0001111000011110", "0001001110110001", "0001000001101001", "0001000000000000", "0001000010000100", "0001001011110110", "0001000001001110", "0001000000000000", "0000111100001111",
 -- Row 12 
 "0100011100011100", "0011001100110011", "0010001000100010", "0001010111001001", "0001000110100111", "0001000100010001", "0001000100011111", "0001001110110001", "0001000100010001", "0001000100010001", "0001000010000100",
 -- Row 13 
 "0100011000100011", "0011001110110111", "0010011101100010", "0001100011111001", "0001001101010010", "0001001001001001", "0001001000100111", "0001010001010001", "0001001001001001", "0001001001001001", "0001000101101010",
 -- Row 14 
 "0100010001000100", "0011010111100101", "0010110010000101", "0001111000011110", "0001010011100101", "0001010000000000", "0001011101000101", "0001010010100101", "0001001110110001", "0001001011110110", "0001001001001001",
 -- Row 15 
 "0011110000111100", "0011100011100011", "0011001100110011", "0010000000000000", "0001100001100001", "0001011001000010", "0001011101000101", "0001010101010101", "0001010010100101", "0001001110110001", "0001001011110110"
);

signal r_a2 : flat_lut :=(
 -- Row 0 
 "0000010110110110", "0000010101110110", "0000111000011111", "0000101100110011", "0000101000110000", "0000101001010010", "0000101011110010", "0000101000100101", "0000100001110100", "0000100101001111", "0000100100011010",
 -- Row 1 
 "0000010110111010", "0000011000000000", "0001001000110100", "0000110101011111", "0000101111111010", "0000110001001100", "0000110110001101", "0000110100000000", "0000101011000010", "0000101111101010", "0000101110110011",
 -- Row 2 
 "0000011001101000", "0000011011100010", "0001100011010011", "0001000101111001", "0000111100110010", "0000111111110100", "0001001001011011", "0001010101000111", "0000111111100011", "0001000101010110", "0001000111001111",
 -- Row 3 
 "0000011011110001", "0000011101110101", "0010011001110101", "0001010101101010", "0001000111001111", "0001001110010011", "0001100110111000", "0001101000110110", "0001010110001110", "0001011011111110", "0001101000000001",
 -- Row 4 
 "0000011101010111", "0000011111000111", "0011011010011101", "0001100101110101", "0001010111001001", "0001100010100011", "0010010000001100", "0010100001110100", "0010011111110110", "0010010000011011", "0011100101111100",
 -- Row 5 
 "0000100000000000", "0000100000011110", "0100010100100001", "0001101101010100", "0001011001001010", "0001100111000010", "0010101011110010", "0010011010001100", "0010101010001110", "0010001010101100", "0011101110010100",
 -- Row 6 
 "0000100011100101", "0000100011110111", "0101000111101011", "0001101101001110", "0001011011101010", "0001101101010100", "0011000100110011", "0010101100011101", "0011011111000110", "0010100010010100", "0100010101011001",
 -- Row 7 
 "0000101000001010", "0000101000100000", "0110010111000011", "0001110111010111", "0001100001100001", "0001110110000101", "0011100101111100", "0010100110011100", "0011100000000011", "0010100011110101", "0100001000110010",
 -- Row 8 
 "0000101110010111", "0000101100100100", "0110000100111100", "0001110101011100", "0001100011010011", "0001110110000101", "0011100011111100", "0010111101111101", "0101000011101000", "0011000100101110", "0101111011111010",
 -- Row 9 
 "0000110010110011", "0000110000110111", "0110011101101000", "0001110110111000", "0001100100011111", "0001111000000001", "0011101001110110", "0010111110101001", "0101101111111010", "0011010000000011", "0110111110001100",
 -- Row 10 
 "0000111000001110", "0000110110000111", "0110111001111000", "0001111001011010", "0001100101110000", "0001111010000110", "0011110010101110", "0010111011001111", "0100101000001101", "0010111011010110", "0100001010011010",
 -- Row 11 
 "0000111101000110", "0000111010110101", "0111011010011110", "0001111100000111", "0001101001111010", "0010000100011011", "0100000001000000", "0011000010001011", "0101010111110010", "0011001100101000", "0100101001001101",
 -- Row 12 
 "0001000011000111", "0001000000101001", "0111101100110111", "0001111111000001", "0001100110011100", "0010000000010000", "0100001101010001", "0011000110111110", "0100011100110100", "0010111010001001", "0100000010111010",
 -- Row 13 
 "0001000111101111", "0001000101000111", "1000000000100000", "0010000011000100", "0001100100111110", "0001111101100011", "0100010011010111", "0011001110000101", "0100110001010100", "0010111101001000", "0100001110100001",
 -- Row 14 
 "0001001010010101", "0001000111101000", "1000000000001100", "0010000100001000", "0001100111100111", "0001111110101000", "0100010011010111", "0011001100110011", "0100101011101010", "0010111000111011", "0100001001010100",
 -- Row 15 
 "0001010000001010", "0001001101010000", "1000001000010001", "0010000011111001", "0001100111001100", "0010000000011101", "0100011001001101", "0011001110110100", "0100110001100001", "0010110111110101", "0100001011010110"
);
 -- Total elements: 176 (16 rows x 11 columns)
signal r_c2 : flat_lut :=(
 -- Row 0 
 "1011011000001011", "1010001111010111", "1000110100111101", "0111111000000111", "0111101001000100", "0111011010111001", "0111000000111000", "0101011000111011", "0100000110001001", "0100101001111001", "0100010001000100",
 -- Row 1 
 "1001110110001001", "1001110110001001", "1000100010001000", "0111010100000111", "0111000111000111", "0110111010110011", "0110100100000110", "0100111000000100", "0011100001111111", "0100000110001001", "0011101010000011",
 -- Row 2 
 "1001010011110010", "1001001001001001", "0111110000011111", "0110110100111010", "0110101001100011", "0110011110110010", "0110000001100000", "0100101001111001", "0011000110100110", "0011110010101110", "0011001100110011",
 -- Row 3 
 "1000101011011000", "1000011001001011", "0111001101100001", "0101101100000101", "0101100100001011", "0101100000010110", "0101001110010111", "0100000110001001", "0010101100011101", "0011011010011101", "0010110110000010",
 -- Row 4 
 "1000010000100001", "0111111000000111", "0110110100111010", "0101001010111111", "0101011100100110", "0101011000111011", "0101000100011011", "0011110010101110", "0010011111110110", "0011000110100110", "0010101100011101",
 -- Row 5 
 "1000001000001000", "0111011010111001", "0110011110110010", "0100101100100111", "0100111000000100", "0100110101001000", "0100101100100111", "0011000000110000", "0010010100111100", "0010110110000010", "0010100011110101",
 -- Row 6 
 "1000000100000010", "0111010100000111", "0110011001100110", "0100010001000100", "0100101001111001", "0100101100100111", "0100100111001101", "0010101100011101", "0010001011011100", "0010101100011101", "0010011100000010",
 -- Row 7 
 "1000000000000000", "0111010000110010", "0110010111000011", "0100001100100101", "0100100100100100", "0100100111001101", "0100011111011100", "0010011100000010", "0001111110000001", "0010100011110101", "0010010100111100",
 -- Row 8 
 "0111111110000000", "0110111001010100", "0110000100111100", "0100001000010000", "0100101001111001", "0100100111001101", "0100011100111100", "0010001110011110", "0001111001010111", "0010011111110110", "0010001110011110",
 -- Row 9 
 "0111111100000001", "0110110111110101", "0110000011110010", "0100000100000100", "0100100111001101", "0100100100100100", "0100010101101100", "0010000011000100", "0001110010111110", "0010011100000010", "0010001011011100",
 -- Row 10 
 "0111111010000100", "0110110110010111", "0110000010101001", "0100000010000001", "0100100100100100", "0100100001111110", "0100010001000100", "0001110101000001", "0001101111000100", "0010011010100100", "0010001000100010",
 -- Row 11 
 "0111111000000111", "0110110100111010", "0110000001100000", "0100000000000000", "0100101001111001", "0100110010001111", "0100010001000100", "0001101101001110", "0001101011011011", "0010011100000010", "0010000101101111",
 -- Row 12 
 "0111110111010110", "0110110100010100", "0110000001000011", "0100000010000001", "0100011100111100", "0100100100100100", "0100010101101100", "0001101001101101", "0001101001000001", "0010011000011010", "0010000011000100",
 -- Row 13 
 "0111110110001100", "0110110011011101", "0110000000011000", "0100000110001001", "0100010101101100", "0100011010011110", "0100010011010111", "0001100111000010", "0001100111000010", "0010010100111100", "0010000000100000",
 -- Row 14 
 "0111110101110011", "0110110011001010", "0110000000001001", "0100001000010000", "0100011100111100", "0100011100111100", "0100010011010111", "0001100110011001", "0001100101001000", "0010010001101000", "0001111110000001",
 -- Row 15 
 "0111110101000010", "0110110010100101", "0101111111101100", "0100000110001001", "0100011010011110", "0100011111011100", "0100010101101100", "0001100100110100", "0001100011010011", "0010001110011110", "0001111011101001"
);

--     --- Debugging signals

    signal r_R0_00 : unsigned(15 downto 0) := "0111111100000000"; -- Debugging signal for R0 value
    signal r_R0_01 : unsigned(15 downto 0) := "0011001000000000"; -- Debugging signal for R0 value

    signal r_R0_21 : unsigned(15 downto 0) := "0000100000000000"; -- Debugging signal for R0 value
    signal r_R0_22 : unsigned(15 downto 0) := "0111101100000000"; -- Debugging signal for R0 value
    signal r_R0_26 : unsigned(15 downto 0) := "0000111100000000"; -- Debugging signal for R0 value
    signal r_R0_55 : unsigned(15 downto 0) := "0101111100000000";

    signal r_c1_00 : unsigned(15 downto 0) := "0100111011000100"; -- Debugging signal for C1 value

    signal dbg_tbl_name : integer range 0 to 5 := 0; -- Debugging signal for table name
begin

  -- Map the internal signal to the entity's output
  o_data <= unsigned(mem_out);

 -- Process for reading and writing data in GHDL with the Flat LUT
process(i_clk)
begin
    if rising_edge(i_clk) then
        if table_name = "R0" then
            dbg_tbl_name <= 1; -- Debugging signal for table name
            r_R0_00 <= r_R0tbl(0); -- Debugging signal for R0 value
            r_R0_01 <= r_R0tbl(1); -- Debugging signal for R0 value
            r_R0_26 <= r_R0tbl(26); -- Debugging signal for R0 value
            r_R0_21 <= r_R0tbl(21); -- Debugging signal for R0 value
            r_R0_55 <= r_R0tbl(55); -- Debugging signal for
            -- Write operation: Store data in the flat LUT at the specified write addresss
            if i_wr_en = '1' then
                if i_waddr < to_unsigned(176, 8) then
                    r_R0tbl(to_integer(i_waddr)) <= i_data; 
                else
                    null;
                end if;
            end if;
            -- Read operation: Output data from the flat LUT at the specified read address
            if i_raddr < to_unsigned(176, 8) then
                mem_out <= std_logic_vector(r_R0tbl(to_integer(i_raddr)));
            else
                mem_out <= std_logic_vector(r_R0tbl(175)); -- Return the last valid entry
            end if;
        elsif table_name = "a1" then
            dbg_tbl_name <= 2; -- Debugging signal for table name
            if i_wr_en = '1' then
                if i_waddr < to_unsigned(176, 8) then
                    r_a1(to_integer(i_waddr)) <= i_data; 
                else
                    null;
                end if;
            end if;
            if i_raddr < to_unsigned(176, 8) then
                mem_out <= std_logic_vector(r_a1(to_integer(i_raddr)));
            else
                mem_out <= std_logic_vector(r_a1(175)); -- Return the last valid entry
            end if;
        elsif table_name = "c1" then
            r_c1_00 <= r_c1(0); -- Debugging signal for C1 value
            dbg_tbl_name <= 3; -- Debugging signal for table name
            if i_wr_en = '1' then
                if i_waddr < to_unsigned(176, 8) then
                    r_c1(to_integer(i_waddr)) <= i_data; 
                else
                    null;
                end if;
            end if;
            if i_raddr < to_unsigned(176, 8) then
                mem_out <= std_logic_vector(r_c1(to_integer(i_raddr)));
            else
                mem_out <= std_logic_vector(r_c1(175)); -- Return the last valid entry
            end if;


        elsif table_name = "a2" then
            dbg_tbl_name <= 4; -- Debugging signal for table name
            if i_wr_en = '1' then
                if i_waddr < to_unsigned(176, 8) then
                    r_a2(to_integer(i_waddr)) <= i_data; 
                else
                    null;
                end if;
            end if;
            if i_raddr < to_unsigned(176, 8) then
                mem_out <= std_logic_vector(r_a2(to_integer(i_raddr)));
            else
                mem_out <= std_logic_vector(r_a2(175)); -- Return the last valid entry
            end if;
        elsif table_name = "c2" then
            dbg_tbl_name <= 5; -- Debugging signal for table name
            if i_wr_en = '1' then
                if i_waddr < to_unsigned(176, 8) then
                    r_c2(to_integer(i_waddr)) <= i_data; 
                else
                    null;
                end if;
            end if;
            if i_raddr < to_unsigned(176, 8) then
                mem_out <= std_logic_vector(r_c2(to_integer(i_raddr)));
            else
                mem_out <= std_logic_vector(r_c2(175)); -- Return the last valid entry
            end if;
        end if;
    end if;
end process;

end architecture rtl;

